module uart_rx #(parameter CLK_FREQ = 100_000_000, parameter BAUD_RATE = 9600) (
    input clk,
    input rx,
    output reg [7:0] data_out,
    output reg rx_done
);
    localparam WAIT_COUNT = CLK_FREQ / BAUD_RATE;
    reg [31:0] count = 0;
    reg [3:0] bit_idx = 0;
    reg [1:0] state = 0;

    always @(posedge clk) begin
        rx_done <= 0;
        case (state)
            0: begin // Idle: Wait for start bit (0)
                count <= 0;
                bit_idx <= 0;
                if (rx == 0) state <= 1;
            end
            1: begin // Start bit: Wait half period to sample in middle
                if (count == WAIT_COUNT / 2) begin
                    count <= 0;
                    state <= 2;
                end else count <= count + 1;
            end
            2: begin // Data bits
                if (count == WAIT_COUNT) begin
                    count <= 0;
                    data_out[bit_idx] <= rx;
                    if (bit_idx == 7) state <= 3;
                    else bit_idx <= bit_idx + 1;
                end else count <= count + 1;
            end
            3: begin // Stop bit
                if (count == WAIT_COUNT) begin
                    rx_done <= 1;
                    state <= 0;
                end else count <= count + 1;
            end
        endcase
    end
endmodule